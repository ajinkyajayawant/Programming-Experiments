module hello_world;

initial begin
$display("Hello world by ajinkya");
#10$finish;
end

endmodule
