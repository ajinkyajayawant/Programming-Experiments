module DFlipFlop(d,clk,Q,qB);
	input d,clk;
	
